`timescale 1ns / 1ps
`include "defines.v"
module prv32_ALU(
    input   wire [31:0] a, b,
    input   wire [4:0]  shamt,
    output  reg  [31:0] r,
    output  wire        cf, zf, vf, sf,
    input   wire [4:0]  alufn
);
    wire [31:0] add, sub, op_b;
    wire cfa, cfs;
    
    assign op_b = (~b);
    assign {cf, add} = alufn[0] ? (a + op_b + 1'b1) : (a + b);
    
    assign zf = (add == 0);
    assign sf = add[31];
    assign vf = (a[31] ^ (op_b[31]) ^ add[31] ^ cf);
    
    wire[31:0] sh;
    shifter shifter0(a, shamt, alufn[1:0], sh);
    reg[63:0]m,ms,msu;

    always @ * begin
        r = 0;
        (* parallel_case *)
        case (alufn)
            `ALU_ADD: r = add;
            `ALU_SUB : r = add;
            `ALU_PASS : r = b;
            `ALU_OR:  r = a | b;
            `ALU_AND:  r = a & b;
            `ALU_XOR:  r = a ^ b;
            `ALU_SRL:  r=sh;
            `ALU_SLL:  r=sh;
            `ALU_SRA:  r=sh;
            `ALU_SLT:  r = {31'b0,(sf != vf)}; 
            `ALU_SLTU:  r = {31'b0,(~cf)};  
            
            `ALU_MUL :  begin ms=$signed(a) *$signed(b); r=ms[31:0]; end
            `ALU_MULHU: begin m = a*b; r=m[63:32]; end
            `ALU_MULH:  begin ms=$signed(a) *$signed(b); r=ms[63:32]; end
            `ALU_MULHSU: begin msu= $signed(a)* b; r=msu[63:32]; end
            
            // ★★★ 나눗셈(DIV, REM) 완전 제거 ★★★
            // 여기 있던 코드들을 다 지웠습니다. 주석 처리도 불안하니 그냥 없앱니다.
            
            default: r = 32'b0;
        endcase
    end
endmodule